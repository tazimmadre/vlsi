`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "interface.sv"
`include "environment.sv"
`include "tbench_top.sv"
`include "test.sv"
`include "design.sv"